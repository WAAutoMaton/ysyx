import "DPI-C" function void difftest_signal_up(
    input int pc,
    input int regs_0, input int regs_1, input int regs_2, input int regs_3,
    input int regs_4, input int regs_5, input int regs_6, input int regs_7,
    input int regs_8, input int regs_9, input int regs_10, input int regs_11,
    input int regs_12, input int regs_13, input int regs_14, input int regs_15,
    input int regs_16, input int regs_17, input int regs_18, input int regs_19,
    input int regs_20, input int regs_21, input int regs_22, input int regs_23,
    input int regs_24, input int regs_25, input int regs_26, input int regs_27,
    input int regs_28, input int regs_29, input int regs_30, input int regs_31,
    input int csr_0, input int csr_1, input int csr_2, input int csr_3, input int csr_4, input int csr_5
);
module DiffTestSignal(
  input         enable,
  input  [31:0] pc,
  input  [31:0] regs_0,
  input  [31:0] regs_1,
  input  [31:0] regs_2,
  input  [31:0] regs_3,
  input  [31:0] regs_4,
  input  [31:0] regs_5,
  input  [31:0] regs_6,
  input  [31:0] regs_7,
  input  [31:0] regs_8,
  input  [31:0] regs_9,
  input  [31:0] regs_10,
  input  [31:0] regs_11,
  input  [31:0] regs_12,
  input  [31:0] regs_13,
  input  [31:0] regs_14,
  input  [31:0] regs_15,
  input  [31:0] regs_16,
  input  [31:0] regs_17,
  input  [31:0] regs_18,
  input  [31:0] regs_19,
  input  [31:0] regs_20,
  input  [31:0] regs_21,
  input  [31:0] regs_22,
  input  [31:0] regs_23,
  input  [31:0] regs_24,
  input  [31:0] regs_25,
  input  [31:0] regs_26,
  input  [31:0] regs_27,
  input  [31:0] regs_28,
  input  [31:0] regs_29,
  input  [31:0] regs_30,
  input  [31:0] regs_31,
  input  [31:0] csr_0,
  input  [31:0] csr_1,
  input  [31:0] csr_2,
  input  [31:0] csr_3,
  input  [31:0] csr_4,
  input  [31:0] csr_5
);
	always @(*) begin
	  if (enable) begin 
	  	difftest_signal_up(
			pc,
			regs_0,
			regs_1,
			regs_2,
			regs_3,
			regs_4,
			regs_5,
			regs_6,
			regs_7,
			regs_8,
			regs_9,
			regs_10,
			regs_11,
			regs_12,
			regs_13,
			regs_14,
			regs_15,
			regs_16,
			regs_17,
			regs_18,
			regs_19,
			regs_20,
			regs_21,
			regs_22,
			regs_23,
			regs_24,
			regs_25,
			regs_26,
			regs_27,
			regs_28,
			regs_29,
			regs_30,
			regs_31,
			csr_0,
			csr_1,
			csr_2,
			csr_3,
			csr_4,
			csr_5
		);
	  end
	end
endmodule
